module mul2 (input logic [31:0] d0,
             output logic [31:0] y);

    always_comb
    begin
        y = d0;
    end

endmodule
